							-------------------------------------------------------------------------------------------------
							-------------------------------------------------------------------------------------------------
							-------------------------------------------------------------------------------------------------
							----  *   )                                                                                  ----
							----` )  /( (      )      (    (           (  (  (            (    (   (   (          (  (   ----
							---- ( )(_)))\    (      ))\   )\    (     )\))( )\   (      ))\  ))\  )(  )\   (     )\))(  ----
							----(_(_())((_)   )\  ' /((_) ((_)   )\ ) ((_))\((_)  )\ )  /((_)/((_)(()\((_)  )\ ) ((_))\  ----
							----|_   _| (_) _((_)) (_))   | __| _(_/(  (()(_)(_) _(_/( (_)) (_))   ((_)(_) _(_/(  (()(_) ----
							----  | |   | || '  \()/ -_)  | _| | ' \))/ _` | | || ' \))/ -_)/ -_) | '_|| || ' \))/ _` |  ----
							----  |_|   |_||_|_|_| \___|  |___||_||_| \__, | |_||_||_| \___|\___| |_|  |_||_||_| \__, |  ----
							----                                      |___/                                      |___/   ----
							-------------------------------------------------------------------------------------------------
							-------------------------------------------------------------------------------------------------
							-------------------------------------------------------------------------------------------------

------------------------------------------------------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------------------------------------------------------
----           _____     _                      ___             __ _     _                                       _              __ _  ----
----    o O O |_   _|   (_)    _ __     ___    | __|   _ _     / _` |   (_)    _ _      ___     ___      _ _    (_)    _ _     / _` | ----
----   o        | |     | |   | '  \   / -_)   | _|   | ' \    \__, |   | |   | ' \    / -_)   / -_)    | '_|   | |   | ' \    \__, | ----
----  TS__[O]  _|_|_   _|_|_  |_|_|_|  \___|   |___|  |_||_|   |___/   _|_|_  |_||_|   \___|   \___|   _|_|_   _|_|_  |_||_|   |___/  ----
---- {======|_|"""""|_|"""""|_|"""""|_|"""""|_|"""""|_|"""""|_|"""""|_|"""""|_|"""""|_|"""""|_|"""""|_|"""""|_|"""""|_|"""""|_|"""""| ----
----./o--000'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-'"`-0-0-' ----
------------------------------------------------------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------------------------------------------------------

-------------------------------------DESCRIPTION------------------------------------------
------------------------------------------------------------------------------------------
-- Bridge da FIFO 8bit to AXI4 Stream.													--
------------------------------------------------------------------------------------------
------------------------------------------------------------------------------------------


library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	
entity AXI4Stream_RS232_v1_0_M00_AXIS_RX is
	generic (
		-- Width of S_AXIS address bus. The slave accepts the read and write addresses of width C_M_AXIS_TDATA_WIDTH.
		C_M_AXIS_TDATA_WIDTH	: integer	:= 8
	);
	port (
		--------------FIFO_DATA (8bit)--------------
		--FIFO_DATA_rst 				: OUT 	STD_LOGIC; Reset lo da chi scrive la FIFO
		FIFO_DATA_clk 				: OUT 	STD_LOGIC;
		FIFO_DATA_dout 				: IN 	STD_LOGIC_VECTOR(8-1 DOWNTO 0);
		FIFO_DATA_rd_en 			: OUT 	STD_LOGIC;
		FIFO_DATA_empty				: IN 	STD_LOGIC;
		FIFO_DATA_almost_empty 		: IN 	STD_LOGIC;
		--------------------------------------------
		
		----------------AXI4-Stream-----------------
		-- AXI4Stream Clock
		M_AXIS_ACLK		: IN 	STD_LOGIC;
		-- AXI4Stream Reset
		M_AXIS_ARESETN	: IN 	STD_LOGIC;
		-- Master Stream Ports. TVALID indicates that the master is driving a valid transfer, A transfer takes place when both TVALID and TREADY are asserted. 
		M_AXIS_TVALID	: OUT 	STD_LOGIC;
		-- TDATA is the primary payload that is used to provide the data that is passing across the interface from the master.
		M_AXIS_TDATA	: OUT 	STD_LOGIC_VECTOR(C_M_AXIS_TDATA_WIDTH-1 DOWNTO 0);
		-- TREADY indicates that the slave can accept a transfer in the current cycle.
		M_AXIS_TREADY	: IN 	STD_LOGIC
		--------------------------------------------
	);
end AXI4Stream_RS232_v1_0_M00_AXIS_RX;

architecture implementation of AXI4Stream_RS232_v1_0_M00_AXIS_RX is
	
	----------------------------SIGNALS-----------------------------
	signal M_AXIS_TVALID_int	: STD_LOGIC;
	----------------------------------------------------------------

begin
	
	---------DIRECT ASSIGNMENT----------
	FIFO_DATA_clk			<= M_AXIS_ACLK;
	--FIFO_DATA_rst 			<= not M_AXIS_ARESETN;
	
	M_AXIS_TDATA			<= FIFO_DATA_dout;
	
	FIFO_DATA_rd_en			<= M_AXIS_TREADY and M_AXIS_TVALID_int;
	
	M_AXIS_TVALID_int		<= not FIFO_DATA_empty and M_AXIS_ARESETN;
	M_AXIS_TVALID			<= M_AXIS_TVALID_int;

	------------------------------------

end implementation;